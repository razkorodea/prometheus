-------------------------------------------------------------------------------
-- SIAE MICROELETTRONICA
-------------------------------------------------------------------------------
--   FILENAME :   thesis.vhd
--
--     AUTHOR :   Gheorghe Balan        
-- START DATE :   xx/yy/zzzz
-------------------------------------------------------------------------------
-- DESCRIPTION 
--		> ...
-------------------------------------------------------------------------------
-- NOTES 
--		> ...
-------------------------------------------------------------------------------
-- CHANGES 
-- 	> ...
--
--
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ============================================================================
-- ENTITY
-- ============================================================================

entity thesis is
end thesis;


-- ============================================================================
-- ARCHITECTURE
-- ============================================================================

architecture rtl of thesis is

   ----------------------------------------------------------------------------
   -- CONSTANTS
   ----------------------------------------------------------------------------


   ----------------------------------------------------------------------------
   -- COMPONENTS
   ----------------------------------------------------------------------------


   ----------------------------------------------------------------------------
   -- NETS
   ----------------------------------------------------------------------------


begin

end rtl;