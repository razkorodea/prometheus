-------------------------------------------------------------------------------
-- SIAE MICROELETTRONICA
-------------------------------------------------------------------------------
--   FILENAME :   krypto_pkg.vhd
-- 
--     AUTHOR :   Gheorghe Balan        
-- START DATE :   xx/yy/zzzz
-------------------------------------------------------------------------------
-- DESCRIPTION 
--		> ...
-------------------------------------------------------------------------------
-- NOTES 
--		> ...
-------------------------------------------------------------------------------
-- CHANGES 
-- 	> ...
-- 
-- 
--

 
library ieee;
use ieee.std_logic_1164.all;



package krypto_pkg is
   ----------------------------------------------------------------------------
   -- 
   ----------------------------------------------------------------------------
   type class_krypto_ctrl is record
      ph_ctrl        : std_logic_vector (31 downto 0);
      ph_init        : std_logic_vector (31 downto 0);
   end record;
   

   
end krypto_pkg;
